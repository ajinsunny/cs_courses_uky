`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:28:59 02/09/2015 
// Design Name: 
// Module Name:    Lab3 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Lab3(
    input [1:0] HAND,
    input GO1,
    input GO2,
    output [2:0] AN,
    output [7:0] SSEG,
    output DISPLAY
    );

endmodule
